module module_antirebote (

//antirebote

//entradas de teclado

//registro de antirebote

//buffer con registro de desplazamiento

 
);
    
endmodule
